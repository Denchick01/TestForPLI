module TestForPLI;
endmodule
