`include "input_driver.v"
`include "time_handler.v"

module TestForPLI;
endmodule
